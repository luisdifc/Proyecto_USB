module Registers_Module (CLK);
//outputs declaration


//inputs declaration
input wire CLK;


endmodule