module Reset_Module (CLK);
//outputs declaration


//inputs declaration
input wire CLK;

//STATE MACHINE
always @(posedge CLK) begin 
	
end //always @(posedge CLK)

endmodule