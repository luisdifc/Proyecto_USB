module Registros(ADDR, RNW, WR_DATA, RD_DATA, req, ACK);

input [7:0] ADDR, RD_DATA, WR_DATA;
input RNW, req, ACK;

reg [15:0] VENDOR_ID, PRODUCT_ID, DEVICE_ID, USBTYPEC_REV, USBPD_REV_VER, PD_INTERFACE_REV, ALERT, ALERT_MASK, DEVICE_CAPABILITIES_1,
		   DEVICE_CAPABILITIES_2, VBUS_VOLTAGE, VBUS_SINK_DISCONNECT_THRESHOLD, VBUS_STOP_DISCHARGE_THRESHOLD, VBUS_VOLTAGE_ALARM_HI_CFG, VBUS_VOLTAGE_ALARM_LO_CFG;

reg [3:0] POWER_STATUS_MASK, FAULT_STATUS_MASK, CONFIG_STANDARD_OUTPUT, TCPC_CONTROL, ROLE_CONTROL, FAULT_CONTROL, POWER_CONTROL, CC_STATUS, POWER_STATUS,
		  FAULT_STATUS, COMMAND, STANDARD_INPUT_CAPABILITIES, STANDARD_OUTPUT_CAPABILITIES, MESSAGE_HEADER_INFO, RECEIVE_DETECT, RECEIVE_BYTE_COUNT, RX_BUF_FRAME_TYPE,
		  RX_BUF_HEADER_BYTE_0, RX_BUF_HEADER_BYTE_1, RX_BUF_OBJ1_BYTE_0, RX_BUF_OBJ1_BYTE_1, RX_BUF_OBJ1_BYTE_2, RX_BUF_OBJ1_BYTE_3, RX_BUF_OBJ2_BYTE_0, RX_BUF_OBJ2_BYTE_1,
		  RX_BUF_OBJ2_BYTE_2, RX_BUF_OBJ2_BYTE_3, RX_BUF_OBJ3_BYTE_0, RX_BUF_OBJ3_BYTE_1, RX_BUF_OBJ3_BYTE_2, RX_BUF_OBJ3_BYTE_3, RX_BUF_OBJ4_BYTE_0, RX_BUF_OBJ4_BYTE_1,
		  RX_BUF_OBJ4_BYTE_2, RX_BUF_OBJ4_BYTE_3, RX_BUF_OBJ5_BYTE_0, RX_BUF_OBJ5_BYTE_1, RX_BUF_OBJ5_BYTE_2, RX_BUF_OBJ5_BYTE_3, RX_BUF_OBJ6_BYTE_0, RX_BUF_OBJ6_BYTE_1,
		  RX_BUF_OBJ6_BYTE_2, RX_BUF_OBJ6_BYTE_3, RX_BUF_OBJ7_BYTE_0, RX_BUF_OBJ7_BYTE_1, RX_BUF_OBJ7_BYTE_2, RX_BUF_OBJ7_BYTE_3, TRANSMIT, TRANSMIT_BYTE_COUNT, 
		  TX_BUF_OBJ1_BYTE_0, TX_BUF_OBJ1_BYTE_1, TX_BUF_OBJ1_BYTE_2, TX_BUF_OBJ1_BYTE_3, TX_BUF_OBJ2_BYTE_0, TX_BUF_OBJ2_BYTE_1, TX_BUF_OBJ2_BYTE_2, TX_BUF_OBJ2_BYTE_3,
		  TX_BUF_OBJ3_BYTE_0, TX_BUF_OBJ3_BYTE_1, TX_BUF_OBJ3_BYTE_2, TX_BUF_OBJ3_BYTE_3, TX_BUF_OBJ4_BYTE_0, TX_BUF_OBJ4_BYTE_1, TX_BUF_OBJ4_BYTE_2, TX_BUF_OBJ4_BYTE_3,
		  TX_BUF_OBJ5_BYTE_0, TX_BUF_OBJ5_BYTE_1, TX_BUF_OBJ5_BYTE_2, TX_BUF_OBJ5_BYTE_3, TX_BUF_OBJ6_BYTE_0, TX_BUF_OBJ6_BYTE_1, TX_BUF_OBJ6_BYTE_2, TX_BUF_OBJ6_BYTE_3,
		  TX_BUF_OBJ7_BYTE_0, TX_BUF_OBJ7_BYTE_1, TX_BUF_OBJ7_BYTE_2, TX_BUF_OBJ7_BYTE_3; 
		  

endmodule
